* File name: C:\Users\Hammad\Desktop\IC Project\SRAM.sch
* Software version: DSCH 3.5
* Created 16/01/2022 17:47:38
*
* Voltage and current sources
*
VBTN1 2 0 DC 0 PULSE(0 1.0 1.00N 0.1N 0.1N 1.00N 3.00N )
VBTN2 3 0 DC 0 PULSE(0 1.0 2.00N 0.1N 0.1N 2.00N 5.00N )
vdd 1 0 DC 1.0
VBTN3 6 0 DC 0 PULSE(0 1.0 3.00N 0.1N 0.1N 3.00N 7.00N )
*
* Passive devices
*
*
* Active devices
*
MN1 3 2 4 3 MN W=0.3u L=0.07u
MP1 4 5 1 4 MP W=0.5u L=0.07u
MN2 4 5 0 4 MN W=0.3u L=0.07u
MN3 0 4 5 0 MN W=0.3u L=0.07u
MP2 1 4 5 1 MP W=0.5u L=0.07u
MN4 5 2 6 5 MN W=0.3u L=0.07u
*
* Warning: "spice.lib" not found, model not declared
.TRAN 0.1ns 250ns
* Dump time and volts in "SRAM.txt"
.control
run
set nobreak
print  V(2) V(3) V(6)  V(5) V(4)  > SRAM.txt
plot  V(2) V(3) V(6)  V(5) V(4) 
.endc
.OPTIONS DELMIN=0 RELTOL=1E-6
.END
